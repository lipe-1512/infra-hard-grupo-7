module and_branch (
    input in1,
    output out
);
    assign out = 1'b1 && in1;
    
endmodule